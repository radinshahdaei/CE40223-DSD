
`include "little_endian_mem.v"

module little_endian_mem_tb();

    reg [15:0] addr;
    reg [1:0] byte_sel;
    reg we, re, clk;
    reg [31:0] data;

    wire [31:0] read_data;
    wire [7:0] data_out_byte;

    little_endian_mem uut (
        .addr(addr),
        .byte_sel(byte_sel),
        .we(we),
        .re(re),
        .clk(clk),
        .data(data),
        .read_data(read_data),
        .data_out_byte(data_out_byte)
    );

    initial begin
        clk = 0;
        forever #5 clk = !clk;
    end

    initial begin
        addr = 0;
        byte_sel = 0;
        we = 0;
        re = 0;
        data = 0;
addr = 16'hFBE1;
data = 32'h13482835;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1FD7;
data = 32'hDBC262ED;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h691F;
data = 32'h8582180D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1E59;
data = 32'h0FF097F6;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA459;
data = 32'h28D516D5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD463;
data = 32'hA7057262;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h69CB;
data = 32'h7B413108;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h46D5;
data = 32'h4FA52BEF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD284;
data = 32'h2D2ACD27;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h26B9;
data = 32'hC5787346;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6BA8;
data = 32'h9E7C3642;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h39D5;
data = 32'h22227BF7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC7B0;
data = 32'h3A9512A9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0F67;
data = 32'h3D9B6B96;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE52F;
data = 32'hF1F76C7F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD308;
data = 32'h1677E787;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5A49;
data = 32'h0929BCEB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAF28;
data = 32'hE1B4CC23;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2457;
data = 32'h395C191B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAE82;
data = 32'hB11647E6;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9759;
data = 32'hFE58E29B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4DC1;
data = 32'h322E4176;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8BDF;
data = 32'h2E982BA8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0E14;
data = 32'hD8513000;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h796A;
data = 32'h9F8F51D7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF1E9;
data = 32'hA360EE70;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6CCB;
data = 32'hF9DF32D5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD8D2;
data = 32'hB2AF15C8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6EE0;
data = 32'h8C424A83;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB020;
data = 32'hC23736DB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h557E;
data = 32'h263FDA4D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFE5A;
data = 32'h563EF079;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFA53;
data = 32'h35B719D7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB1C5;
data = 32'hE04599E8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h229C;
data = 32'hA1A3E0EE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAB3D;
data = 32'hF7138BC9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3D20;
data = 32'h9CC0EADD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3FC2;
data = 32'h885C994A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF56F;
data = 32'hAD4065B4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB99F;
data = 32'h484D61EF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF1E1;
data = 32'hA6611A89;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6122;
data = 32'hA710D199;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDDD4;
data = 32'hC94393F4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEB17;
data = 32'h9E4B6EFF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0F92;
data = 32'hC9134A6B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2B35;
data = 32'h4AADC5EC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC86C;
data = 32'hA49406D8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCCAD;
data = 32'h52260E22;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0589;
data = 32'h01279A33;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5B7F;
data = 32'h7ADE7498;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB689;
data = 32'h8B1CC89E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEB1E;
data = 32'hA3BD4403;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB2E6;
data = 32'h1A617CD7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h904E;
data = 32'h86302EB6;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEB92;
data = 32'hF99051E0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDC8D;
data = 32'hA0D9E2BA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCAAA;
data = 32'hE66ADF98;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB9D8;
data = 32'h361680A0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h01B7;
data = 32'h5C49780C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5329;
data = 32'h445043A0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0294;
data = 32'h7D4A8077;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4403;
data = 32'h8514A454;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h89AD;
data = 32'h3860C2A7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC6D1;
data = 32'h67D6718E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE4FE;
data = 32'h1892B515;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0956;
data = 32'h7247BD2A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6935;
data = 32'hBCEEAA00;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBAA4;
data = 32'h5524D6C8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE205;
data = 32'h626793E1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h438D;
data = 32'hE8D8EDB6;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hACCE;
data = 32'hC2D2704D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA57A;
data = 32'h17BC4EA7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB5DC;
data = 32'hED1309C9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3FA7;
data = 32'hD9C03ED5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE10B;
data = 32'h8BE8EBD4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD211;
data = 32'hAF23E3CE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8977;
data = 32'hF2C78EFF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8BEF;
data = 32'hBB186C76;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC437;
data = 32'h267575B4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC8F2;
data = 32'h7B323549;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFDC2;
data = 32'hFC43E7AE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7BE9;
data = 32'hCA8E7C29;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5283;
data = 32'hB7F1C275;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB3C0;
data = 32'h82B47E76;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h235F;
data = 32'hBBEE66BE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBB09;
data = 32'hC4E3E42C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB62B;
data = 32'h7EAD37D5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0C01;
data = 32'h022778F0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB009;
data = 32'h46988D24;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3F31;
data = 32'hAF4411BE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFDE1;
data = 32'hB7FF19F9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDCDE;
data = 32'h5AA2B754;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h95E5;
data = 32'hDE06BF30;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h90D7;
data = 32'hDE7F5F1D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5965;
data = 32'h31A9B201;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4CA3;
data = 32'hD03C82F3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h49B2;
data = 32'hD9471C69;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4345;
data = 32'hC83A5807;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8237;
data = 32'h366754A5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0E8E;
data = 32'h813A480A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h76C4;
data = 32'hD27F5A99;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEA04;
data = 32'h77D88C83;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8A00;
data = 32'hF72AC9BC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4719;
data = 32'hA3A772F1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h09D0;
data = 32'h63C512AF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h041E;
data = 32'h6CB7712D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h65C8;
data = 32'h5761FE8E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4CB9;
data = 32'hD43BF008;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h17AF;
data = 32'hF8522A71;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h25C0;
data = 32'h31A59ADC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h996B;
data = 32'h9A908C88;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5798;
data = 32'hAC45D2F7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h97E7;
data = 32'h016FB666;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h60F0;
data = 32'h0960B551;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h192F;
data = 32'h8BA8E5EA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDD07;
data = 32'hB6B191DF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEC33;
data = 32'h59E14A86;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2B77;
data = 32'hAEE6DC25;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h01A1;
data = 32'h53003B3D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1971;
data = 32'h0F497180;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD1E3;
data = 32'h4B98C842;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5967;
data = 32'hBB47AF1D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC812;
data = 32'hD8EBE2BC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5B28;
data = 32'h04A0A231;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAED1;
data = 32'hE2BC9C96;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF3E5;
data = 32'h0210BA44;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCCCF;
data = 32'h5063C5CC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7638;
data = 32'h8228C583;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC866;
data = 32'h0BDEB458;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2C1B;
data = 32'hAA5A75E5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB369;
data = 32'h552DCC00;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE217;
data = 32'h8722A265;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7D3C;
data = 32'h3B3E1F50;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h73FC;
data = 32'hB5477B02;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h33CE;
data = 32'hC933F124;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA580;
data = 32'h2BED4695;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4611;
data = 32'hF0B957F7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5920;
data = 32'hBB49FA67;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDCB8;
data = 32'h829595D1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6307;
data = 32'h1FFE1931;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8A1F;
data = 32'hCA0246CA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h52C7;
data = 32'h35AD5785;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFC33;
data = 32'h6A11D0F0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3728;
data = 32'hF4898CA3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA1FC;
data = 32'hCC9EB4C8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC631;
data = 32'h909740AF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h32CA;
data = 32'h8A5A20DF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4F64;
data = 32'hBE4ECAE8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h39E5;
data = 32'hA8E74890;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBF13;
data = 32'h0C03B245;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD756;
data = 32'hC33DB765;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h729E;
data = 32'h3F4C578D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEE6C;
data = 32'h36612D18;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9B22;
data = 32'h4BDE3836;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB120;
data = 32'h7A251E8D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8F4C;
data = 32'h8521E143;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5208;
data = 32'h8A2FA12F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1360;
data = 32'h1DAE07E7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h639B;
data = 32'hE2E66490;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h656B;
data = 32'hF80FCEE0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4C19;
data = 32'h1D6A729C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h07C7;
data = 32'hAB609B7B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAA9E;
data = 32'hBE795F92;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC81C;
data = 32'hDD5E4FE2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF3A6;
data = 32'hCE0DAEA4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFBAE;
data = 32'h3934CDCC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h097D;
data = 32'h862BD959;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1A30;
data = 32'hF1082F14;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE9C8;
data = 32'h8FBDF054;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6955;
data = 32'hBACBFCB2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFFC7;
data = 32'h5E110CE9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3B82;
data = 32'h74DD26DB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h106F;
data = 32'h1F8CE5B9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC5AF;
data = 32'h6AB4589F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA64A;
data = 32'hE9A8CD22;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h621D;
data = 32'h337BC101;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5A98;
data = 32'hE6D502F6;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6180;
data = 32'h117CECE8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8C2B;
data = 32'h6D9ED996;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0900;
data = 32'h95A643C9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB415;
data = 32'hF9C7BF88;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAA38;
data = 32'h9213BAF2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEA68;
data = 32'hD07C3664;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h93E6;
data = 32'h56CAF62C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h786C;
data = 32'hBED4E8BE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8F84;
data = 32'hB5E497CE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4B55;
data = 32'hC81483F9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6AB2;
data = 32'h4093AB4C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA6B3;
data = 32'h01960486;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h30CF;
data = 32'h8E6F6DBF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h41CE;
data = 32'h2F2B38FE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5DD8;
data = 32'h9E652845;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8F9F;
data = 32'h931AC731;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4C00;
data = 32'h9051679B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h00D2;
data = 32'hE05F94D4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB162;
data = 32'h7417B08A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h879B;
data = 32'h688AF5A1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h713D;
data = 32'h0CB03113;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h030A;
data = 32'h499BF814;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h028F;
data = 32'h781B06F2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3005;
data = 32'h535D83E5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5CC8;
data = 32'h777107FC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD5EF;
data = 32'h4D51FC1B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBD5A;
data = 32'hC04EE610;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h598B;
data = 32'hE79EC396;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0E58;
data = 32'hBCC063AA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h085D;
data = 32'h013E73E6;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0287;
data = 32'h6F7A7AF2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF8C2;
data = 32'h593CD403;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6C3A;
data = 32'h4BED4E96;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB313;
data = 32'h3BEE7B83;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC4B8;
data = 32'h83F3D859;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h936B;
data = 32'h67B528CA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6FB6;
data = 32'h23E3C9BB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0433;
data = 32'hA78CBF74;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC8F0;
data = 32'hC3398223;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9735;
data = 32'h20EE1266;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6F49;
data = 32'h6F38CD0B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h07AB;
data = 32'hEB8D7A2B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h73D9;
data = 32'hDBC322BF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA1A8;
data = 32'hF6E1E4A8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFF91;
data = 32'hAF2204E1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h233B;
data = 32'h4DC486D2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h60D1;
data = 32'hB8DA9D8F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0701;
data = 32'h82E42B76;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6673;
data = 32'hE779E129;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3EE1;
data = 32'hE61BFF7D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC0F0;
data = 32'hC71623DD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE1B8;
data = 32'h7D50A719;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA63C;
data = 32'h3BBD5CED;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAE38;
data = 32'h6B3CCAFA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFF98;
data = 32'hF698579F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0422;
data = 32'hAFA465BD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0D00;
data = 32'h93F757D4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2545;
data = 32'h6ADCB60B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8416;
data = 32'h986CFC4B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h20B0;
data = 32'h49C0EFDB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h328E;
data = 32'h00C53A2B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h580B;
data = 32'h5C64DC1A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA57D;
data = 32'h03D827D1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h28D2;
data = 32'h6685041E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB477;
data = 32'h37E786FA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1ABB;
data = 32'h02BF87EB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1580;
data = 32'h4B9F746B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC9EC;
data = 32'hC531B06C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAC89;
data = 32'hAC0631E9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h968A;
data = 32'hE096D156;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2207;
data = 32'h81065577;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFF77;
data = 32'hFC3F1970;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h15E1;
data = 32'hD75CAB62;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h554E;
data = 32'hC009B153;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC21D;
data = 32'hEFFA1F9E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h85CA;
data = 32'h904AE971;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB22E;
data = 32'h9F1E83F4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF0FE;
data = 32'h7ED263D1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAF36;
data = 32'h625FDB9F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5C3B;
data = 32'hEBFB2617;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3BD1;
data = 32'h3ADCDE6C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h66BB;
data = 32'h75813AE5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF7C3;
data = 32'hE64EC44E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8030;
data = 32'h784CB3C1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h377E;
data = 32'hC1DA6D82;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDC12;
data = 32'h8A4CD496;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1212;
data = 32'h36518C4B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF1A1;
data = 32'h3990AB2F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h33F6;
data = 32'h3CCE11AD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5CB7;
data = 32'h183B83FC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC999;
data = 32'h78E87ECC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4CD8;
data = 32'h34D988A4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h58B0;
data = 32'h53E5CE7B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD89F;
data = 32'h4D8C15D4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h387F;
data = 32'hB5C38058;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC36D;
data = 32'h8EEBF096;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDC90;
data = 32'h222DE483;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8F33;
data = 32'hF9ED68E1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3409;
data = 32'h011C060A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9004;
data = 32'h259FE53E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD6F5;
data = 32'h9B5D45F5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE35D;
data = 32'h3A30A332;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3AA8;
data = 32'h9530DE78;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE900;
data = 32'h88A81CB2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h547E;
data = 32'h087149BF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h22E2;
data = 32'h8633E11E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3221;
data = 32'h4226FF93;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFF19;
data = 32'h64781A0B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5230;
data = 32'hFE677BC3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE03D;
data = 32'h4190B8EA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6905;
data = 32'h24CFACDE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h89BF;
data = 32'hB7DC3A10;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA31B;
data = 32'hF4CCC502;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD154;
data = 32'h1F2E20E3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2C12;
data = 32'h9519C13E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h277E;
data = 32'h8C69DA9C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5512;
data = 32'h45F1BE54;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h01EB;
data = 32'h3987E033;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h83C3;
data = 32'hB8E90CC9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4B09;
data = 32'h67C4DAC9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0DF7;
data = 32'h3D72F3B3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h43B9;
data = 32'h5C7B7552;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCE25;
data = 32'hBB894B49;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3F45;
data = 32'h34B336B3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1742;
data = 32'hE6E1525F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE395;
data = 32'h7B48D9B0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC333;
data = 32'h541D9868;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hED53;
data = 32'h0399717C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h43D0;
data = 32'hE753922F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h752E;
data = 32'h5124AF51;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2A06;
data = 32'hBBC699AC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCF3E;
data = 32'hCA994624;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDEDA;
data = 32'h56C4B0D8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0A56;
data = 32'h3C9CA8EC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h143D;
data = 32'hACC04B66;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9747;
data = 32'hFC286BE3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h227F;
data = 32'h85F42E70;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE0D3;
data = 32'hA0FE38FF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB59F;
data = 32'h61A1BC21;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9AE1;
data = 32'h008A5F63;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD35F;
data = 32'h6324E026;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9C11;
data = 32'hA19B887A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h42BB;
data = 32'h28AEE773;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7BC2;
data = 32'h16A176A7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h64D9;
data = 32'h94E16FF1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h19C6;
data = 32'hE31309AC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6027;
data = 32'h71D696BE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC080;
data = 32'h04BB1523;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3CE3;
data = 32'hC8651DE1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h201E;
data = 32'h120E8532;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h74F5;
data = 32'hD514D2FE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9128;
data = 32'h1CA43E3E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC354;
data = 32'hE5473BE2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2786;
data = 32'h6E255C16;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h625B;
data = 32'h8B36B691;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA082;
data = 32'hA1E2490D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEA92;
data = 32'hD918D789;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1E34;
data = 32'hD5711620;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4314;
data = 32'h215C7C99;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8606;
data = 32'hB6F52B3D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5A93;
data = 32'h9EC86AE6;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD41C;
data = 32'h8970DA2E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6357;
data = 32'hE7BB7476;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4E13;
data = 32'hA0EACC6D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h895C;
data = 32'h5009C308;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h16DF;
data = 32'h656A7D7D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3D04;
data = 32'hFF9611CF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3311;
data = 32'h401E30A4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5390;
data = 32'h70B7FDAC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8A2F;
data = 32'h9D5F6F26;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB34F;
data = 32'hA690F12C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2987;
data = 32'h83AC3370;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB599;
data = 32'h1E15FD2F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCDB9;
data = 32'hAEC6E535;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCFF4;
data = 32'hE828B245;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h635B;
data = 32'h31C5B31A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9FBD;
data = 32'hF684FFFF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4417;
data = 32'h9392B82A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h629D;
data = 32'h86F23DB4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h362F;
data = 32'hA65C986F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA762;
data = 32'hAD34C832;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h954C;
data = 32'h9611F312;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1F26;
data = 32'hB3943B2E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC446;
data = 32'hD46B24A3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD805;
data = 32'hF45FF3D9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3487;
data = 32'hCDC238F9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5E2E;
data = 32'hC9A9247F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h79B8;
data = 32'hF0C081CD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1F16;
data = 32'h1DF95383;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1189;
data = 32'hBD6FF719;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9A79;
data = 32'h15B78130;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEE6E;
data = 32'hDC862838;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF51D;
data = 32'h8AB19AC4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0CA3;
data = 32'h835A83B4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h513B;
data = 32'h60261558;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3F08;
data = 32'h7EB5B7D9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h23D7;
data = 32'h0B71D80B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hED76;
data = 32'hE05A3387;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBCC6;
data = 32'hCDFD931E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h087F;
data = 32'h8B5A997F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB2AD;
data = 32'hA7D625FB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5B0D;
data = 32'h4B2103B5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF552;
data = 32'hD34C9B19;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hECD5;
data = 32'h0C32B4C6;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFE85;
data = 32'h174EE52A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h45F4;
data = 32'h0530B0BE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h92E1;
data = 32'h7535F2CC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8450;
data = 32'h04D75674;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h33EE;
data = 32'h3CED4651;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCF69;
data = 32'h4DE2699C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5FC1;
data = 32'hE47A6E5A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA3E6;
data = 32'h68B971A2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5C61;
data = 32'hE08F1B92;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h81F9;
data = 32'h442A484B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB1C9;
data = 32'hD5930E40;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB127;
data = 32'h0D6B43F8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB0D1;
data = 32'hF068AF65;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA06B;
data = 32'hD835294E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6DC2;
data = 32'h26946D16;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8207;
data = 32'hA8188BEB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1AE9;
data = 32'h53DCB5EE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8583;
data = 32'h9179262B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE514;
data = 32'h2298275D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2603;
data = 32'hD617416F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD895;
data = 32'h3A79EC61;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h198F;
data = 32'h297A86D1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2D0B;
data = 32'hCC43363F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE618;
data = 32'h182FB863;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF26F;
data = 32'h0B355A32;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFC03;
data = 32'h47276254;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB60D;
data = 32'h1E728FEA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6560;
data = 32'hA07401C8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB731;
data = 32'h7F5EB835;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h19B5;
data = 32'hB13574C0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2222;
data = 32'hD0FBFC16;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEDF3;
data = 32'h382ADD25;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCCE5;
data = 32'h7A45643B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6BD2;
data = 32'h90232841;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF954;
data = 32'h8E477080;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4F4C;
data = 32'hF7B5B691;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h68C4;
data = 32'hF8C53676;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB237;
data = 32'hD99C968B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDF05;
data = 32'h5164554A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE2CF;
data = 32'h768576B3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD849;
data = 32'hB1CAF7BC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5D85;
data = 32'hA59A0AE2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h003F;
data = 32'h1FA4C38C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCBD5;
data = 32'hD35155E7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9E63;
data = 32'h3769BAE3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h40A6;
data = 32'h34D8F11E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7D18;
data = 32'hCFD68B0E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h147C;
data = 32'hE6280FF3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE234;
data = 32'h79CA7128;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9C04;
data = 32'h84705647;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB846;
data = 32'h2388DB0F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA329;
data = 32'h8AE4A094;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5311;
data = 32'h8C3432DD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h78B5;
data = 32'h7656407C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDDBE;
data = 32'hD0C72D0F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4662;
data = 32'hDC0DD801;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h50F1;
data = 32'h0AA4D99B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h79FA;
data = 32'hB6A11E0B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA38A;
data = 32'h2C56FD29;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB573;
data = 32'hC006F305;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5A57;
data = 32'h35D14DDC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3E1A;
data = 32'hBE232A67;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7692;
data = 32'h6AFBA8B3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h33E4;
data = 32'h74C3FBAB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB3C9;
data = 32'h5088957C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCA16;
data = 32'hD2144908;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1CDD;
data = 32'h1594F3EC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7F55;
data = 32'hE2B69F5A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h01C1;
data = 32'h7ED9EB84;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2A81;
data = 32'hD6DD6EE6;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h64FD;
data = 32'h61D0BCD1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0654;
data = 32'h94175D9D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB0CE;
data = 32'h6A02CC75;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8D78;
data = 32'h3B6FB37A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6D73;
data = 32'h53BB7871;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8666;
data = 32'h7BB71A91;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCC48;
data = 32'h6EAA5F14;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7A5D;
data = 32'h87238E83;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8473;
data = 32'hC50CA57C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4C6F;
data = 32'hBD1570A1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h664D;
data = 32'h365DB126;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF44A;
data = 32'h74557D55;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h992A;
data = 32'h6FBDB9E3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE107;
data = 32'h363666CD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE371;
data = 32'h4F780B7D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1C07;
data = 32'hA047A3BC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAEDD;
data = 32'hAE8B16EA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7610;
data = 32'h30931B6D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5D06;
data = 32'hD8AA187A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD6DF;
data = 32'h439AECEB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h615E;
data = 32'h12CA8046;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7059;
data = 32'h41B6F1E7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h31DA;
data = 32'h929F4697;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h32F1;
data = 32'h8456BF38;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8568;
data = 32'h90A86C80;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8A87;
data = 32'h69279E06;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5E42;
data = 32'h60A9BF90;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h07AB;
data = 32'hC8434791;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3EEE;
data = 32'h1F09AB62;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2326;
data = 32'h3904E5B5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6897;
data = 32'h21BD498A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBD05;
data = 32'h7D8EE91F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB447;
data = 32'h7181442F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h577A;
data = 32'hB97A392F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD184;
data = 32'h7F392A23;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4C3C;
data = 32'hE142B0B5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBC13;
data = 32'h1801D768;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDB96;
data = 32'h9F616EED;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB708;
data = 32'h43DAE320;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA670;
data = 32'h87D6FADB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5E66;
data = 32'h667DD7EF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h51FB;
data = 32'hA50236C0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE88C;
data = 32'h2F12841D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8D81;
data = 32'h6AABB695;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h672E;
data = 32'h6F80656A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h53D5;
data = 32'hEBF1C813;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA11B;
data = 32'h449FD626;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h808F;
data = 32'hC050B0D1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6B4E;
data = 32'hFC134BC5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4355;
data = 32'hAFE487AA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB85B;
data = 32'h0F4DED5F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEF19;
data = 32'hBC0E429B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4B35;
data = 32'h81D473C3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB972;
data = 32'hE0FC09E5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2FA6;
data = 32'h5AD6AF40;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h73BA;
data = 32'h495CE280;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5F0A;
data = 32'h05A53EEA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h174D;
data = 32'h724ADD69;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0778;
data = 32'h8A555636;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h01A1;
data = 32'hCDBFBD5F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1AA5;
data = 32'hFD218832;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4917;
data = 32'h4903FDB9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h11D5;
data = 32'hAFAB2004;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE7DE;
data = 32'h272E791C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h04FC;
data = 32'hAF138EB0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h82F4;
data = 32'hACFD5346;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h24D9;
data = 32'h0142CC01;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC15A;
data = 32'h6C99EDDF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC71B;
data = 32'h42D8F946;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h20B8;
data = 32'h5BACC116;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3836;
data = 32'hC4551043;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7409;
data = 32'h0F1CE0AC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF39E;
data = 32'h015FB153;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1D80;
data = 32'hE2012ABD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h543A;
data = 32'hFEAADE65;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h958A;
data = 32'hABA024ED;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7893;
data = 32'h64F4D7CF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE1EA;
data = 32'h543755AC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5504;
data = 32'h217F2201;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h282D;
data = 32'h47D6A794;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6479;
data = 32'hE601D397;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE311;
data = 32'h9B4742FB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA94C;
data = 32'hAC0A42DB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1825;
data = 32'h85C11B7D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6A0E;
data = 32'h818496C8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD58A;
data = 32'hA8562BFE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD9DA;
data = 32'h182CBCDF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA94E;
data = 32'h5B304A41;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0236;
data = 32'hAF04CA9E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF99B;
data = 32'hFC5EF547;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE2F5;
data = 32'h92A16F8C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDF98;
data = 32'hF00AAA5D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5DB5;
data = 32'h9A22E15E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB586;
data = 32'hDA968CC3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h186A;
data = 32'hB78D4BFD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7D26;
data = 32'hF4D2BC09;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3B00;
data = 32'hEE69561A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7715;
data = 32'h05EE9E2C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCBCD;
data = 32'h9017BC00;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3BFF;
data = 32'hB8F39E2E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB8FE;
data = 32'hD3CD60EB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0AE8;
data = 32'h77824471;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h952D;
data = 32'hA772CEDE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9F8C;
data = 32'h97709CCA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h66E0;
data = 32'hD88CC247;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3FB8;
data = 32'hBBF2174B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEE41;
data = 32'hA3F7D23C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9766;
data = 32'h5887CC0D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4881;
data = 32'hC9389370;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBB6B;
data = 32'h03F62A9B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA04E;
data = 32'h2BEFA7BA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1757;
data = 32'hDFB1CF9C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF282;
data = 32'h8DFF8493;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDE79;
data = 32'h3E4EFA1E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA128;
data = 32'hD78140C2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h13A8;
data = 32'h3CBBB6F2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h600A;
data = 32'hD179C576;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0521;
data = 32'hAD27B3DB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7FE8;
data = 32'h98652777;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7551;
data = 32'h8DB58C2A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h20D2;
data = 32'h8F11076F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h66CB;
data = 32'h659FE5BE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4F30;
data = 32'h505ED279;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h53FA;
data = 32'h1E16CBF6;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8C7C;
data = 32'hD13CB614;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCF59;
data = 32'h1A62496D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h87C1;
data = 32'h8FDAD7F1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEAB2;
data = 32'h4637203C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5057;
data = 32'h8E08F8AE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2F62;
data = 32'h34E9941D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDA41;
data = 32'h41643076;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB3D6;
data = 32'h27146FBD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h964A;
data = 32'h49E2C0C3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA103;
data = 32'h755EFB49;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h818E;
data = 32'h4895EF18;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6BEB;
data = 32'h5E939EB4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA09F;
data = 32'h810177E7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8762;
data = 32'h4F06A1E1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFD02;
data = 32'h0009451A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h78E9;
data = 32'h201DAC4C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h682B;
data = 32'hA3FB6E28;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1CA8;
data = 32'hDA3E5B2D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1E8B;
data = 32'h43C573C4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2591;
data = 32'hC792285C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2735;
data = 32'h9153CCF4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3195;
data = 32'hA6EBFF68;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h673C;
data = 32'h41A127BB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB6EB;
data = 32'h5E46C7C4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB746;
data = 32'h44204C25;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1D0D;
data = 32'hB2D3ECA3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7B25;
data = 32'hF6B5A747;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD0DD;
data = 32'h3EF92764;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB808;
data = 32'h32CC1405;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA57C;
data = 32'h1FEB3FF9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3A29;
data = 32'hD46FD518;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCBED;
data = 32'hFAD564B3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2254;
data = 32'h135EE6C1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0691;
data = 32'hFB376593;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDC81;
data = 32'h80B369F2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBA49;
data = 32'h669B8F5D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3ADE;
data = 32'h5A568C52;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h76E1;
data = 32'hA1FC8667;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC871;
data = 32'h58F35153;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1393;
data = 32'h14B6D1BC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0CE2;
data = 32'h112FE3EB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3F46;
data = 32'hAE52C32E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0B34;
data = 32'h68016753;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB6DC;
data = 32'h676F1BC4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB72E;
data = 32'h1E4DC2F1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h18BC;
data = 32'h83AA355C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDD9C;
data = 32'h37D1EA27;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1CF6;
data = 32'hB8E73172;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAE18;
data = 32'hC36ECA5C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC39E;
data = 32'hDCA300B0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9E41;
data = 32'h702B3EC8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFBC3;
data = 32'hD332ADE7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE90C;
data = 32'hCC072656;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB0AB;
data = 32'hACB18A5F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE655;
data = 32'hD255CA1D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h31D3;
data = 32'h177343E7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8C81;
data = 32'hC3469795;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1181;
data = 32'h4EC2E5DB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC3F7;
data = 32'h9DA959F2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCC83;
data = 32'hDE7ACB53;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0E7F;
data = 32'hBF7074C5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBDC8;
data = 32'h878211C2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0135;
data = 32'h65E7993D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB0CD;
data = 32'h9BA384C8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5CF3;
data = 32'hAD674BFA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6B29;
data = 32'h1CF43435;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB07E;
data = 32'hB6A207EA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0974;
data = 32'hBDAD9C68;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD14C;
data = 32'h6F3A8F09;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2BA4;
data = 32'hBEB23CE8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7475;
data = 32'hD8712514;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDE13;
data = 32'h1B75F44C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h626C;
data = 32'h15FFA40C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h283A;
data = 32'h5E781D0E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3BBA;
data = 32'h11AD24C1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h18CD;
data = 32'h92C5CB80;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8588;
data = 32'h6F257B35;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h18C5;
data = 32'hF9325071;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4B86;
data = 32'hBC090F3E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6E9E;
data = 32'h7B32D4C1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4844;
data = 32'h7F015C94;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA945;
data = 32'h32E69B01;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA438;
data = 32'h01A8A499;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2F2A;
data = 32'h0DD0ED62;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9F0C;
data = 32'hE78684F7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5B26;
data = 32'h9C9B0184;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC03F;
data = 32'h86042EA4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h304C;
data = 32'h295AEB5C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6872;
data = 32'hB3BD5E09;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h14C5;
data = 32'h72B005FB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF63B;
data = 32'hBCB10CD9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9DDA;
data = 32'h707AE573;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1A31;
data = 32'h3ECCCE7D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4961;
data = 32'h76644E85;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8E7B;
data = 32'h7A2F721C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h58FF;
data = 32'hE1D3D858;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFB79;
data = 32'h4B179808;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0660;
data = 32'h6388E16B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9E5D;
data = 32'h4460FBBF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4BC1;
data = 32'h6AB0C176;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h33A8;
data = 32'hA43A9958;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE3AE;
data = 32'hA1A36D7E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h698E;
data = 32'h99DA9D1F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h428E;
data = 32'h4CA07C75;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h721C;
data = 32'h90FF9A0F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0859;
data = 32'h82A89789;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAA16;
data = 32'h68DF0E29;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1314;
data = 32'hD2F7A132;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2EF5;
data = 32'h3D0F5A28;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDA87;
data = 32'h2DFBA3AA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8051;
data = 32'h4E934C08;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF6DA;
data = 32'h5528588B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8BBF;
data = 32'h87DB1AFD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h98C2;
data = 32'h9E4FAA75;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1F47;
data = 32'h8CB06C3F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h72DD;
data = 32'hFBE4DD21;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3DB3;
data = 32'h51D632B5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA0A5;
data = 32'h1255CC73;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA7B2;
data = 32'hE2399E90;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h452E;
data = 32'h244AF523;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF589;
data = 32'h19FB3C76;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h951C;
data = 32'h740F6538;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9679;
data = 32'h043EE285;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h18EC;
data = 32'h23149AE6;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h71A3;
data = 32'h2E887408;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4A02;
data = 32'h6FBCFFD1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h938A;
data = 32'hB7C2F485;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hADD7;
data = 32'h0A23AA1E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4E51;
data = 32'h5549FD1C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8624;
data = 32'h1EFCAF17;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC1EB;
data = 32'h11E807CE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h58C0;
data = 32'h1F85C87C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF326;
data = 32'hB89E1729;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF14E;
data = 32'hF6149E62;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCD13;
data = 32'h862ED7A1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2936;
data = 32'h55754B58;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8E52;
data = 32'h734ADDF4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h527B;
data = 32'hFBA80F70;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDD65;
data = 32'hAD11A33B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0A74;
data = 32'h548A627F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC2D7;
data = 32'h47DF7827;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF1B3;
data = 32'hADE3702B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h732B;
data = 32'h1BC3546A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0D69;
data = 32'h1B2E7D16;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h393E;
data = 32'hB05E53A4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1BBF;
data = 32'hBA1039C9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h377B;
data = 32'hE68D29F4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8C7C;
data = 32'hE15A35FB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEDB7;
data = 32'hB386C275;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE2D8;
data = 32'h16772FEB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8BFB;
data = 32'hD1673892;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA28E;
data = 32'h451BCE0E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2627;
data = 32'hFEDA0954;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8BB4;
data = 32'h6066DAE2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2332;
data = 32'h2BB37AAB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2A3A;
data = 32'h658ED759;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h53A0;
data = 32'hE5DBB385;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDF15;
data = 32'h134CB688;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h062B;
data = 32'h7F495A81;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD461;
data = 32'h6AAED8D2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h69D4;
data = 32'hECB95478;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h05F0;
data = 32'hD6EDAF28;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDBE0;
data = 32'hA1CADC7A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFDD4;
data = 32'h3BD2387F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hED8D;
data = 32'h9C148789;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFF22;
data = 32'hBF7979F3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE442;
data = 32'hAEE79872;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9D23;
data = 32'hC3A38D73;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA68D;
data = 32'hB97702CC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4B59;
data = 32'hA2E1441C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD425;
data = 32'h7C9DE366;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h58D8;
data = 32'h072DCC3D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h30A3;
data = 32'hAE599165;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEE58;
data = 32'h8D38F6E4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB34D;
data = 32'hED899BAB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBF42;
data = 32'h98DB87D7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h04ED;
data = 32'hA1A84530;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0A26;
data = 32'hF3653694;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h25CB;
data = 32'hCD479FC9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDB60;
data = 32'h4FCE11A3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h55E4;
data = 32'hFCFDEDC2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF6F7;
data = 32'h3D466DB3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA9C0;
data = 32'h0AAC3165;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3C63;
data = 32'h1B691E0F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h079C;
data = 32'hB356044A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF17D;
data = 32'h62B6C045;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCC86;
data = 32'hC06EF899;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5151;
data = 32'h91313A10;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE95A;
data = 32'hE46B8E81;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC9FB;
data = 32'h760FF7CD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDBB6;
data = 32'hD709A7DF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h73C4;
data = 32'h06A7E6F7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h636A;
data = 32'h08141838;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD4D1;
data = 32'h934AE504;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7CE5;
data = 32'h4F63B976;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h470B;
data = 32'h05775C5D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE3A0;
data = 32'h9EDAA54F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC3CC;
data = 32'h5DD2FC1C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2763;
data = 32'h0055FCE7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h865E;
data = 32'h199F064A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h931D;
data = 32'h26906F32;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAA02;
data = 32'hA87D118B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1B83;
data = 32'h57EB0AD8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFE59;
data = 32'h15B36A5A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD47A;
data = 32'hDDDF2550;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2001;
data = 32'hBCF5B59B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h838F;
data = 32'hF53AC5B1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE1AC;
data = 32'h0ECC1E9F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8315;
data = 32'h90A41C08;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE64B;
data = 32'h7EF1CE85;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4E51;
data = 32'hDBFD7957;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7C79;
data = 32'h6A2EB6D6;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4D1B;
data = 32'h6AD07C24;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA382;
data = 32'hB5BF9AD1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE985;
data = 32'hEAEF0840;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h520E;
data = 32'hB2366B61;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE422;
data = 32'h96000155;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAEB6;
data = 32'hEFAE1F60;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h041D;
data = 32'h35170BFB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCAF0;
data = 32'h737AD541;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6FB1;
data = 32'h3F5B67FD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7021;
data = 32'h3A18B6CB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE153;
data = 32'h86D15D35;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFC4E;
data = 32'hA6C3BCA9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h69DF;
data = 32'hEA5973D1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3289;
data = 32'h3E3D0B72;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9909;
data = 32'hBC053862;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCF0D;
data = 32'hCC2AAFE4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB1F9;
data = 32'h3ACC24DA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE377;
data = 32'hE1E7A1C1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC856;
data = 32'h158E29D5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h46E8;
data = 32'h307D824A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2B35;
data = 32'h7C2BCE26;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4986;
data = 32'h7ECE33A8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h593A;
data = 32'hBD4D736E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1A9A;
data = 32'h2ECBEC8A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2E42;
data = 32'hF83F736C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA4F9;
data = 32'h62E9900C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0861;
data = 32'hCE81DD36;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD063;
data = 32'hEF1FF4F8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h76C6;
data = 32'hDDB1D7BD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h023A;
data = 32'h4FBE6334;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2742;
data = 32'h2EF0D06E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h49E0;
data = 32'hDF735853;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA630;
data = 32'h1228534D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCA18;
data = 32'hD3A239D0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3C72;
data = 32'hE47AB65C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h86F3;
data = 32'h78A87A8B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBDC9;
data = 32'h92A58AA3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h47C4;
data = 32'hD044AD6B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB2F7;
data = 32'h19A8AA69;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0BEE;
data = 32'hDCB186AF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h49F8;
data = 32'h7D21C668;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF7D4;
data = 32'h2E42B0E2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFDDC;
data = 32'h35D6E6A9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1CF3;
data = 32'hD064966D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFFDC;
data = 32'h093B4C09;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB872;
data = 32'hF8F866C0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAC84;
data = 32'hC2F4CC5B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3B65;
data = 32'hFED13C1A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF7A3;
data = 32'h9663B1CA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF3DD;
data = 32'h3869A064;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB56A;
data = 32'h966E084E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6220;
data = 32'hF71DDA27;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4EE6;
data = 32'h52465148;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1794;
data = 32'hF216BD04;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC490;
data = 32'hF2507662;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9A85;
data = 32'h013C9FF8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBF26;
data = 32'h57B9C269;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9352;
data = 32'h2408602A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7803;
data = 32'h29538F57;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h648E;
data = 32'hFCF68CFD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE62A;
data = 32'h881176E0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h98AA;
data = 32'hEFE8BAD7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC79E;
data = 32'hAE8CA9F2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8FBF;
data = 32'hC05A586C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8F65;
data = 32'h2574D844;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF783;
data = 32'h350DEC13;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3CA8;
data = 32'h69822557;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBB22;
data = 32'h9761E41B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD93E;
data = 32'h7F05929D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h30EB;
data = 32'hF86CCDC1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5DEA;
data = 32'hC9453E23;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDD0E;
data = 32'h873C6DE1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8EB4;
data = 32'h7C19EBD4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCE7E;
data = 32'hE4DE9F09;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h96C3;
data = 32'h9860F319;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9B5D;
data = 32'h854B32B4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDC6A;
data = 32'h5CD2BBCA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1726;
data = 32'hFAB8325E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9B06;
data = 32'h86583A08;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h851A;
data = 32'hACE242BC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE6F3;
data = 32'h99D4B07A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h35AE;
data = 32'h8F5AD552;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9059;
data = 32'h3FC14163;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h06E2;
data = 32'hF6686C27;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9679;
data = 32'h49053E19;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h43DF;
data = 32'hFF1EB47C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h323B;
data = 32'h42840ECE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h37D9;
data = 32'h8492E932;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1BD2;
data = 32'h314E5E41;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF344;
data = 32'hEBAC0389;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h59D9;
data = 32'h0568D2DC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7B08;
data = 32'hC9EF08DE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCF64;
data = 32'hCAC45109;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDCAF;
data = 32'h54FB7F3E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB422;
data = 32'hEA2F0479;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4F6F;
data = 32'hEB238E96;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB4F9;
data = 32'hA1D50C44;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h089D;
data = 32'hF8B8A0BE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8123;
data = 32'h737B5D13;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5510;
data = 32'h8AD357C1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9F2C;
data = 32'h50B72976;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB5CA;
data = 32'h1258F0D9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBB3D;
data = 32'hF8C03E43;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCE7A;
data = 32'hF6297969;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1580;
data = 32'hC2516003;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h80A0;
data = 32'h84F923B4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h32CE;
data = 32'h508A3C38;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE74D;
data = 32'hF73FD60A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h180E;
data = 32'hBE1EDC40;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9FCE;
data = 32'hB1BD2FDB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3B75;
data = 32'h684C77D0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h20FE;
data = 32'hC021DF01;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5FA1;
data = 32'h4FA88912;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h39E7;
data = 32'h969FF0A8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0EB6;
data = 32'h474795FC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9B0A;
data = 32'hA35ABB7F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF563;
data = 32'hBC18AADA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE730;
data = 32'h5A5BDF11;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE524;
data = 32'hB6E4142F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEA99;
data = 32'h897E3F9E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h36FA;
data = 32'h3ED5EF24;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4C60;
data = 32'h2F1DA551;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h48FE;
data = 32'hA4FCF916;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4367;
data = 32'h9AFF9CC7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD880;
data = 32'h1577F88E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC887;
data = 32'h55C44E4A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD937;
data = 32'h9047B039;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFC70;
data = 32'h5B1423FF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4935;
data = 32'hE3D5CEE2;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h38AD;
data = 32'hF6615DE1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA16E;
data = 32'hD4708C03;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h650E;
data = 32'h2307F90A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2959;
data = 32'h0D240449;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h56B6;
data = 32'hAF1B2EFD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h226F;
data = 32'h9CC44BBC;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h99E9;
data = 32'hC8BE2195;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE95F;
data = 32'hC5E147F0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0CF1;
data = 32'h254165B3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hCB7A;
data = 32'h4161EE33;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2DA9;
data = 32'hCDABE934;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDEF5;
data = 32'h98B95A24;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h80A1;
data = 32'hFFCFB8F0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC259;
data = 32'h83A981BE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3E5E;
data = 32'h98A91FC3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h13C2;
data = 32'h15002A09;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h32A0;
data = 32'h9000B4EA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h65FD;
data = 32'h4E99CDA3;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3666;
data = 32'h81A133D8;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h923B;
data = 32'h2E45DB86;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5758;
data = 32'h3A2B6C05;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3AC1;
data = 32'hE479A096;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF6F8;
data = 32'h091E4404;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD3DA;
data = 32'h9A7FC49D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD679;
data = 32'h0F447246;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h1F1C;
data = 32'h2A43177C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3847;
data = 32'hC6758960;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC3C1;
data = 32'h2372B879;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEB62;
data = 32'h5307848B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB7DF;
data = 32'h975DA3B1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h72B4;
data = 32'hBB9E93DA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h2072;
data = 32'h4706B903;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE6EC;
data = 32'hFF2961D1;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3DF9;
data = 32'h8FDA7ED5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4F10;
data = 32'hD17DE2C9;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEFE1;
data = 32'hF8EEC5CA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8105;
data = 32'h1D697466;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8798;
data = 32'hD2217AA7;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h6ADB;
data = 32'h713E7AC0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h89EE;
data = 32'hC3FC154B;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8801;
data = 32'h22C0B942;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h51FE;
data = 32'hCD6BED6F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD6E7;
data = 32'h52279AFB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hBC06;
data = 32'h03B9B974;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h743E;
data = 32'hAE270CA4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEA0D;
data = 32'h670B0A3C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hD352;
data = 32'hE28664CD;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4FF0;
data = 32'h7C467AE5;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h4109;
data = 32'h9F8EAE5F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h5DBF;
data = 32'hCD3D0665;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h3763;
data = 32'h8C4E1323;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hEDEA;
data = 32'h1B35BA37;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA4F3;
data = 32'h9F7EFCEF;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC9CC;
data = 32'h8FFB4EC6;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7720;
data = 32'hFFEF7A41;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h09CA;
data = 32'hC277D458;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h632A;
data = 32'h80674461;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h27C6;
data = 32'h3C2EB74C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h692B;
data = 32'hE016B76D;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h556B;
data = 32'h918ED589;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAA1C;
data = 32'hE282171F;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h27C3;
data = 32'h355D6967;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF268;
data = 32'h73BC961E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA62C;
data = 32'hE68C9C24;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hAD85;
data = 32'h1470030C;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hDA0E;
data = 32'hA1053A20;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h79CF;
data = 32'h0A5B1D57;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h30CE;
data = 32'h8A1A9E47;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hE041;
data = 32'hDF22A316;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h0A00;
data = 32'h05392BAE;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hC2B8;
data = 32'h76EBF472;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h44C1;
data = 32'h8085761A;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h73B8;
data = 32'hD9E75588;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7B4D;
data = 32'hDF6B43CB;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h9FD3;
data = 32'h2585AE4E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hF8D5;
data = 32'h7252FDDA;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h17A1;
data = 32'hC22C2AB6;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hA764;
data = 32'hD2695D16;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hB035;
data = 32'hDECF6E60;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hADE5;
data = 32'h7EF993D4;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8C46;
data = 32'hE8E845E0;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8DC6;
data = 32'hA3A2E369;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h7699;
data = 32'hE111C639;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'h8E1E;
data = 32'h83EB3B9E;
we = 1;
#10;
we = 0;
$display("Written %h to address %h", data, addr);
#10;
addr = 16'hFBE1;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1FD7;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h691F;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1E59;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA459;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD463;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h69CB;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h46D5;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD284;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h26B9;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6BA8;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h39D5;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC7B0;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0F67;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE52F;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD308;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5A49;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAF28;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2457;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAE82;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9759;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4DC1;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8BDF;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0E14;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h796A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF1E9;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6CCB;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD8D2;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6EE0;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB020;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h557E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFE5A;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFA53;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB1C5;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h229C;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAB3D;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3D20;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3FC2;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF56F;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB99F;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF1E1;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6122;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDDD4;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEB17;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0F92;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2B35;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC86C;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCCAD;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0589;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5B7F;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB689;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEB1E;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB2E6;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h904E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEB92;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDC8D;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCAAA;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB9D8;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h01B7;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5329;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0294;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4403;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h89AD;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC6D1;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE4FE;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0956;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6935;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBAA4;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE205;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h438D;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hACCE;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA57A;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB5DC;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3FA7;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE10B;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD211;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8977;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8BEF;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC437;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC8F2;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFDC2;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7BE9;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5283;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB3C0;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h235F;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBB09;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB62B;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0C01;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB009;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3F31;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFDE1;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDCDE;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h95E5;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h90D7;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5965;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4CA3;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h49B2;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4345;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8237;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0E8E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h76C4;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEA04;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8A00;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4719;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h09D0;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h041E;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h65C8;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4CB9;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h17AF;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h25C0;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h996B;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5798;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h97E7;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h60F0;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h192F;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDD07;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEC33;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2B77;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h01A1;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1971;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD1E3;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5967;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC812;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5B28;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAED1;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF3E5;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCCCF;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7638;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC866;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2C1B;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB369;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE217;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7D3C;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h73FC;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h33CE;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA580;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4611;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5920;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDCB8;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6307;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8A1F;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h52C7;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFC33;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3728;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA1FC;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC631;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h32CA;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4F64;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h39E5;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBF13;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD756;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h729E;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEE6C;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9B22;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB120;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8F4C;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5208;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1360;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h639B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h656B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4C19;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h07C7;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAA9E;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC81C;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF3A6;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFBAE;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h097D;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1A30;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE9C8;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6955;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFFC7;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3B82;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h106F;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC5AF;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA64A;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h621D;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5A98;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6180;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8C2B;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0900;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB415;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAA38;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEA68;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h93E6;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h786C;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8F84;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4B55;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6AB2;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA6B3;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h30CF;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h41CE;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5DD8;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8F9F;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4C00;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h00D2;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB162;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h879B;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h713D;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h030A;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h028F;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3005;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5CC8;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD5EF;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBD5A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h598B;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0E58;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h085D;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0287;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF8C2;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6C3A;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB313;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC4B8;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h936B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6FB6;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0433;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC8F0;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9735;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6F49;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h07AB;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h73D9;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA1A8;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFF91;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h233B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h60D1;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0701;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6673;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3EE1;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC0F0;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE1B8;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA63C;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAE38;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFF98;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0422;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0D00;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2545;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8416;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h20B0;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h328E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h580B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA57D;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h28D2;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB477;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1ABB;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1580;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC9EC;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAC89;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h968A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2207;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFF77;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h15E1;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h554E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC21D;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h85CA;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB22E;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF0FE;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAF36;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5C3B;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3BD1;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h66BB;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF7C3;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8030;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h377E;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDC12;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1212;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF1A1;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h33F6;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5CB7;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC999;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4CD8;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h58B0;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD89F;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h387F;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC36D;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDC90;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8F33;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3409;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9004;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD6F5;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE35D;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3AA8;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE900;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h547E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h22E2;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3221;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFF19;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5230;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE03D;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6905;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h89BF;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA31B;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD154;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2C12;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h277E;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5512;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h01EB;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h83C3;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4B09;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0DF7;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h43B9;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCE25;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3F45;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1742;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE395;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC333;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hED53;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h43D0;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h752E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2A06;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCF3E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDEDA;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0A56;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h143D;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9747;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h227F;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE0D3;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB59F;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9AE1;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD35F;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9C11;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h42BB;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7BC2;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h64D9;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h19C6;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6027;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC080;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3CE3;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h201E;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h74F5;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9128;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC354;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2786;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h625B;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA082;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEA92;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1E34;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4314;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8606;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5A93;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD41C;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6357;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4E13;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h895C;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h16DF;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3D04;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3311;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5390;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8A2F;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB34F;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2987;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB599;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCDB9;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCFF4;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h635B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9FBD;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4417;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h629D;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h362F;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA762;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h954C;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1F26;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC446;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD805;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3487;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5E2E;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h79B8;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1F16;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1189;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9A79;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEE6E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF51D;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0CA3;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h513B;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3F08;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h23D7;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hED76;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBCC6;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h087F;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB2AD;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5B0D;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF552;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hECD5;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFE85;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h45F4;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h92E1;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8450;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h33EE;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCF69;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5FC1;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA3E6;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5C61;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h81F9;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB1C9;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB127;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB0D1;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA06B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6DC2;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8207;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1AE9;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8583;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE514;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2603;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD895;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h198F;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2D0B;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE618;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF26F;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFC03;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB60D;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6560;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB731;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h19B5;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2222;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEDF3;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCCE5;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6BD2;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF954;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4F4C;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h68C4;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB237;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDF05;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE2CF;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD849;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5D85;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h003F;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCBD5;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9E63;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h40A6;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7D18;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h147C;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE234;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9C04;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB846;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA329;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5311;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h78B5;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDDBE;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4662;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h50F1;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h79FA;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA38A;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB573;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5A57;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3E1A;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7692;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h33E4;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB3C9;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCA16;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1CDD;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7F55;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h01C1;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2A81;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h64FD;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0654;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB0CE;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8D78;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6D73;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8666;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCC48;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7A5D;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8473;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4C6F;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h664D;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF44A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h992A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE107;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE371;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1C07;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAEDD;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7610;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5D06;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD6DF;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h615E;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7059;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h31DA;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h32F1;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8568;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8A87;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5E42;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h07AB;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3EEE;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2326;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6897;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBD05;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB447;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h577A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD184;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4C3C;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBC13;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDB96;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB708;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA670;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5E66;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h51FB;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE88C;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8D81;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h672E;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h53D5;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA11B;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h808F;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6B4E;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4355;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB85B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEF19;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4B35;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB972;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2FA6;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h73BA;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5F0A;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h174D;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0778;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h01A1;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1AA5;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4917;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h11D5;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE7DE;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h04FC;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h82F4;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h24D9;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC15A;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC71B;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h20B8;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3836;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7409;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF39E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1D80;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h543A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h958A;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7893;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE1EA;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5504;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h282D;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6479;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE311;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA94C;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1825;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6A0E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD58A;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD9DA;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA94E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0236;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF99B;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE2F5;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDF98;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5DB5;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB586;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h186A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7D26;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3B00;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7715;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCBCD;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3BFF;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB8FE;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0AE8;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h952D;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9F8C;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h66E0;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3FB8;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEE41;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9766;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4881;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBB6B;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA04E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1757;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF282;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDE79;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA128;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h13A8;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h600A;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0521;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7FE8;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7551;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h20D2;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h66CB;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4F30;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h53FA;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8C7C;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCF59;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h87C1;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEAB2;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5057;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2F62;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDA41;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB3D6;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h964A;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA103;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h818E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6BEB;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA09F;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8762;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFD02;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h78E9;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h682B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1CA8;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1E8B;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2591;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2735;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3195;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h673C;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB6EB;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB746;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1D0D;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7B25;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD0DD;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB808;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA57C;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3A29;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCBED;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2254;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0691;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDC81;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBA49;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3ADE;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h76E1;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC871;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1393;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0CE2;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3F46;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0B34;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB6DC;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB72E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h18BC;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDD9C;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1CF6;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAE18;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC39E;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9E41;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFBC3;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE90C;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB0AB;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE655;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h31D3;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8C81;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1181;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC3F7;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCC83;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0E7F;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBDC8;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0135;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB0CD;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5CF3;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6B29;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB07E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0974;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD14C;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2BA4;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7475;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDE13;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h626C;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h283A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3BBA;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h18CD;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8588;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h18C5;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4B86;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6E9E;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4844;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA945;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA438;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2F2A;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9F0C;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5B26;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC03F;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h304C;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6872;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h14C5;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF63B;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9DDA;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1A31;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4961;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8E7B;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h58FF;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFB79;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0660;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9E5D;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4BC1;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h33A8;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE3AE;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h698E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h428E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h721C;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0859;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAA16;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1314;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2EF5;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDA87;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8051;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF6DA;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8BBF;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h98C2;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1F47;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h72DD;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3DB3;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA0A5;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA7B2;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h452E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF589;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h951C;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9679;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h18EC;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h71A3;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4A02;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h938A;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hADD7;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4E51;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8624;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC1EB;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h58C0;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF326;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF14E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCD13;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2936;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8E52;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h527B;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDD65;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0A74;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC2D7;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF1B3;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h732B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0D69;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h393E;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1BBF;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h377B;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8C7C;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEDB7;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE2D8;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8BFB;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA28E;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2627;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8BB4;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2332;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2A3A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h53A0;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDF15;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h062B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD461;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h69D4;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h05F0;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDBE0;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFDD4;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hED8D;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFF22;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE442;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9D23;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA68D;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4B59;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD425;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h58D8;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h30A3;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEE58;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB34D;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBF42;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h04ED;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0A26;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h25CB;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDB60;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h55E4;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF6F7;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA9C0;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3C63;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h079C;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF17D;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCC86;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5151;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE95A;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC9FB;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDBB6;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h73C4;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h636A;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD4D1;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7CE5;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h470B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE3A0;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC3CC;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2763;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h865E;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h931D;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAA02;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1B83;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFE59;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD47A;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2001;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h838F;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE1AC;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8315;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE64B;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4E51;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7C79;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4D1B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA382;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE985;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h520E;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE422;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAEB6;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h041D;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCAF0;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6FB1;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7021;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE153;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFC4E;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h69DF;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3289;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9909;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCF0D;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB1F9;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE377;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC856;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h46E8;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2B35;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4986;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h593A;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1A9A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2E42;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA4F9;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0861;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD063;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h76C6;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h023A;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2742;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h49E0;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA630;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCA18;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3C72;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h86F3;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBDC9;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h47C4;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB2F7;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0BEE;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h49F8;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF7D4;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFDDC;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1CF3;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFFDC;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB872;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAC84;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3B65;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF7A3;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF3DD;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB56A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6220;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4EE6;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1794;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC490;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9A85;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBF26;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9352;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7803;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h648E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE62A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h98AA;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC79E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8FBF;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8F65;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF783;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3CA8;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBB22;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD93E;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h30EB;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5DEA;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDD0E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8EB4;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCE7E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h96C3;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9B5D;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDC6A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1726;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9B06;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h851A;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE6F3;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h35AE;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9059;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h06E2;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9679;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h43DF;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h323B;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h37D9;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1BD2;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF344;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h59D9;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7B08;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCF64;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDCAF;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB422;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4F6F;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB4F9;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h089D;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8123;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5510;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9F2C;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB5CA;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBB3D;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCE7A;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1580;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h80A0;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h32CE;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE74D;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h180E;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9FCE;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3B75;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h20FE;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5FA1;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h39E7;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0EB6;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9B0A;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF563;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE730;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE524;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEA99;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h36FA;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4C60;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h48FE;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4367;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD880;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC887;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD937;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hFC70;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4935;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h38AD;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA16E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h650E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2959;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h56B6;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h226F;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h99E9;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE95F;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0CF1;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hCB7A;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2DA9;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDEF5;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h80A1;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC259;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3E5E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h13C2;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h32A0;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h65FD;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3666;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h923B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5758;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3AC1;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF6F8;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD3DA;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD679;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h1F1C;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3847;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC3C1;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEB62;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB7DF;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h72B4;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h2072;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE6EC;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3DF9;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4F10;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEFE1;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8105;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8798;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h6ADB;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h89EE;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8801;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h51FE;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD6E7;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hBC06;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h743E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEA0D;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hD352;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4FF0;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h4109;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h5DBF;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h3763;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hEDEA;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA4F3;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC9CC;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7720;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h09CA;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h632A;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h27C6;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h692B;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h556B;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAA1C;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h27C3;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF268;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA62C;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hAD85;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hDA0E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h79CF;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h30CE;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hE041;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h0A00;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hC2B8;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h44C1;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h73B8;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7B4D;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h9FD3;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hF8D5;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h17A1;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hA764;
byte_sel = 2'b10;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hB035;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'hADE5;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8C46;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8DC6;
byte_sel = 2'b01;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h7699;
byte_sel = 2'b00;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
addr = 16'h8E1E;
byte_sel = 2'b11;
re = 1;
#10;
$display("Read full data at address %h: %h", addr, read_data);
$display("Byte %h at address %h: %h", byte_sel, addr, data_out_byte);
re = 0;
#10;
        $display("Test completed.");
        $finish;
    end

endmodule
